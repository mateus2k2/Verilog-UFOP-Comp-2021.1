module ex1(A,B);

input A;  //declarar uma entrada;
output B; //declarar uma saida;

assign B=A;

endmodule